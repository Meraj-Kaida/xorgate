module xorgate(a,b,y);

input a,b;//input values
output y;
assign y=a^b;
endmodule
//

